`ifndef XCTCMSG_NETWORKS_SVH
`define XCTCMSG_NETWORKS_SVH

`include "xctcmsg_networks/bus.svh"

`ifdef XCTCMSG_NETWORK_BUS
  `define XCTCMSG_NETWORK_INTERFACE `XCTCMSG_NETWORK_BUS_INTERFACE
  `define XCTCMSG_NETWORK_ADAPTER   `XCTCMSG_NETWORK_BUS_ADAPTER
`endif

`include "xctcmsg_networks/openpiton.svh"

`ifdef XCTCMSG_NETWORK_OPENPITON
  `define XCTCMSG_NETWORK_INTERFACE `XCTCMSG_NETWORK_OPENPITON_INTERFACE
  `define XCTCMSG_NETWORK_ADAPTER   `XCTCMSG_NETWORK_OPENPITON_ADAPTER
`endif

`endif // XCTCMSG_NETWORKS_SVH
